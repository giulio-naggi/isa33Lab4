-- VHDL Entity HAVOC.FPmul_stage2.interface
--
-- Created by
-- Guillermo Marcus, gmarcus@ieee.org
-- using Mentor Graphics FPGA Advantage tools.
--
-- Visit "http://fpga.mty.itesm.mx" for more info.
--
-- 2003-2004. V1.0
--

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY FPmul_stage2 IS
   PORT( 
      A_EXP           : IN     std_logic_vector (7 DOWNTO 0);
      A_SIG           : IN     std_logic_vector (31 DOWNTO 0);
      B_EXP           : IN     std_logic_vector (7 DOWNTO 0);
      B_SIG           : IN     std_logic_vector (31 DOWNTO 0);
      SIGN_out_stage1 : IN     std_logic;
      clk             : IN     std_logic;
      isINF_stage1    : IN     std_logic;
      isNaN_stage1    : IN     std_logic;
      isZ_tab_stage1  : IN     std_logic;
      EXP_in          : OUT    std_logic_vector (7 DOWNTO 0);
      EXP_neg_stage2  : OUT    std_logic;
      EXP_pos_stage2  : OUT    std_logic;
      SIGN_out_stage2 : OUT    std_logic;
      SIG_in          : OUT    std_logic_vector (27 DOWNTO 0);
      isINF_stage2    : OUT    std_logic;
      isNaN_stage2    : OUT    std_logic;
      isZ_tab_stage2  : OUT    std_logic
   );

-- Declarations

END FPmul_stage2 ;

--
-- VHDL Architecture HAVOC.FPmul_stage2.struct
--
-- Created by
-- Guillermo Marcus, gmarcus@ieee.org
-- using Mentor Graphics FPGA Advantage tools.
--
-- Visit "http://fpga.mty.itesm.mx" for more info.
--
-- Copyright 2003-2004. V1.0
--


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ARCHITECTURE struct OF FPmul_stage2 IS

	component dadda_mul is
		port(	A,B : in std_logic_vector(31 downto 0);
				P : out std_logic_vector(63 downto 0));
	end component;

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL EXP_in_int  : std_logic_vector(7 DOWNTO 0);
   SIGNAL EXP_neg_int, EXP_neg_int_0 : std_logic;
   SIGNAL EXP_pos_int, EXP_pos_int_0, EXP_pos_int_1 : std_logic;
   SIGNAL SIG_in_int  : std_logic_vector(27 DOWNTO 0);
   SIGNAL dout        : std_logic;
   SIGNAL dout1       : std_logic_vector(7 DOWNTO 0);
   SIGNAL mw_I4sum, mw_I4sum_0, mw_I4sum_1, mw_I4sum_2       : std_logic_vector(8 DOWNTO 0);
   SIGNAL prod, prod_1, prod_0        : std_logic_vector(63 DOWNTO 0);
   SIGNAL isINF_stage1_2, isNaN_stage1_2, isZ_tab_stage1_2, SIGN_out_stage1_2    : std_logic;
   SIGNAL MUX_EXPR, MUX_EXPR_0    : std_logic;

	component REG is 
	generic (n : integer := 8);
	port(CLK: in std_logic;
		IN_DATA: in std_logic_vector(n-1 downto 0);
		OUT_DATA: out std_logic_vector(n-1 downto 0));
	end component;
	component flipflop is 
		port(CLK: in std_logic;
			IN_DATA: in std_logic;
			OUT_DATA: out std_logic);
	end component;

BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 sig
   -- eb1 1
   SIG_in_int <= prod(47 DOWNTO 20);

   -- HDL Embedded Text Block 2 inv
   -- eb5 5
   EXP_in_int <= (NOT dout1(7)) & dout1(6 DOWNTO 0);

   -- HDL Embedded Text Block 3 latch
   -- eb2 2
   
   PROCESS(clk)
   BEGIN
      IF RISING_EDGE(clk) THEN
         EXP_in <= EXP_in_int;
         SIG_in <= SIG_in_int;
         EXP_pos_stage2 <= EXP_pos_int;
         EXP_neg_stage2 <= EXP_neg_int;
      END IF;
   END PROCESS;

   -- HDL Embedded Text Block 4 latch2
   -- latch2 4
   PROCESS(clk)
   BEGIN
      IF RISING_EDGE(clk) THEN
         isINF_stage2 <= isINF_stage1;
         isNaN_stage2 <= isNaN_stage1;
         isZ_tab_stage2 <= isZ_tab_stage1;
         SIGN_out_stage2 <= SIGN_out_stage1;
      END IF;
   END PROCESS;

   -- HDL Embedded Text Block 5 eb1
   -- exp_pos 5
   EXP_pos_int_0 <= A_EXP(7) AND B_EXP(7);
--   EXP_neg_int <= NOT(A_EXP(7) OR B_EXP(7));
   MUX_EXPR_0 <= '1' WHEN ( (A_EXP(7)='0' AND NOT (A_EXP=X"7F")) AND (B_EXP(7)='0' AND NOT (B_EXP=X"7F")) ) ELSE '0';
   EXP_neg_int_0 <= '1' WHEN MUX_EXPR='1' ELSE '0';


   -- ModuleWare code(v1.1) for instance 'I4' of 'add'
   I4combo: PROCESS (A_EXP, B_EXP)
   VARIABLE mw_I4t0 : std_logic_vector(8 DOWNTO 0);
   VARIABLE mw_I4t1 : std_logic_vector(8 DOWNTO 0);
   VARIABLE mw_I4t01 : unsigned(8 DOWNTO 0);
   BEGIN
      mw_I4t0 := '0' & A_EXP;
      mw_I4t1 := '0' & B_EXP;
	  mw_I4t01 := unsigned(mw_I4t0) + unsigned(mw_I4t1);
      mw_I4sum_0 <= std_logic_vector(mw_I4t01);
   END PROCESS I4combo;
   
   I4combo_1: PROCESS (mw_I4sum_1, dout)
   VARIABLE mw_I4carry : std_logic;
   VARIABLE mw_I4sum_2_0: unsigned(8 DOWNTO 0);
   BEGIN
      mw_I4carry := dout;
	  mw_I4sum_2_0 := unsigned(mw_I4sum_1) + mw_I4carry;
	  mw_I4sum_2 <= std_logic_vector(mw_I4sum_2_0); 
   END PROCESS I4combo_1;
   
   dout1 <= mw_I4sum(7 DOWNTO 0);
   
   -- ModuleWare code(v1.1) for instance 'I2' of 'mult'
   -- I2combo : PROCESS (A_SIG, B_SIG)
   -- VARIABLE dtemp : unsigned(63 DOWNTO 0);
   -- BEGIN
      -- dtemp := (unsigned(A_SIG) * unsigned(B_SIG));
      -- prod_0 <= std_logic_vector(dtemp);
   -- END PROCESS I2combo;
   
   DADDA: dadda_mul port map(A => A_SIG, B => B_SIG, P => prod_0);

	reg_1: reg generic map (n => 64) port map(CLK => clk, IN_DATA => prod_0, OUT_DATA => prod_1);
	reg_2: reg generic map (n => 64) port map(CLK => clk, IN_DATA => prod_1, OUT_DATA => prod);
	reg_3: flipflop port map(CLK => clk, IN_DATA => isINF_stage1, OUT_DATA => isINF_stage1_2);
	reg_4: flipflop port map(CLK => clk, IN_DATA => isINF_stage1_2, OUT_DATA => isINF_stage2);
	reg_5: flipflop port map(CLK => clk, IN_DATA => isNaN_stage1, OUT_DATA => isNaN_stage1_2);
	reg_6: flipflop port map(CLK => clk, IN_DATA => isNaN_stage1_2, OUT_DATA => isINF_stage2);
	reg_7: flipflop port map(CLK => clk, IN_DATA => isZ_tab_stage1, OUT_DATA => isZ_tab_stage1_2);
	reg_8: flipflop port map(CLK => clk, IN_DATA => isZ_tab_stage1_2, OUT_DATA => isZ_tab_stage2);
	reg_9: flipflop port map(CLK => clk, IN_DATA => SIGN_out_stage1, OUT_DATA => SIGN_out_stage1_2);
	reg_10: flipflop port map(CLK => clk, IN_DATA => SIGN_out_stage1_2, OUT_DATA => SIGN_out_stage2);
	reg_11: reg generic map (n => 9) port map(CLK => clk, IN_DATA => mw_I4sum_0, OUT_DATA => mw_I4sum_1);
	reg_12: reg generic map (n => 9) port map(CLK => clk, IN_DATA => mw_I4sum_2, OUT_DATA => mw_I4sum);
	reg_13: flipflop port map(CLK => clk, IN_DATA => MUX_EXPR_0, OUT_DATA => MUX_EXPR);
	reg_14: flipflop port map(CLK => clk, IN_DATA => EXP_neg_int_0, OUT_DATA => EXP_neg_int);
	reg_15: flipflop port map(CLK => clk, IN_DATA => EXP_pos_int_0, OUT_DATA => EXP_pos_int_1);
	reg_16: flipflop port map(CLK => clk, IN_DATA => EXP_pos_int_1, OUT_DATA => EXP_pos_int);
   -- ModuleWare code(v1.1) for instance 'I6' of 'vdd'
   dout <= '1';

   -- Instance port mappings.

END struct;
